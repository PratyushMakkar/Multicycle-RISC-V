`define SIM
`define ICE_40