package rv32I_core_package;

endpackage